module L1_cache(

input clk,
input rst_n,

input lsu_req,
output [DW-1:0] lsu_rdata

);




endmodule

